library ieee;
use ieee.std_logic_1164.all;
use work.all;

entity RSA is
  port(
    -- input
    clk: in std_ulogic;
    -- output
  );
end RSA;
  
  
  
architecture behaviour of RSA is
  -- internal signals
begin -- logic
  -- include RSA_Core
  -- include RSA_Ctrl
end behaviour;
