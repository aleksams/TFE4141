library ieee;
use ieee.std_logic_1164.all;
use work.all;

entity RSA_Ctrl is
  port(
    -- input
    clk: in std_ulogic;
    -- output
  );
end RSA_Ctrl;
  
  
  
architecture behaviour of RSA_Ctrl is
  -- internal signals
begin -- logic

end behaviour;
