library ieee;
use ieee.std_logic_1164.all;
use work.all;

entity RSA_Core is
  port(
    -- input
    clk: in std_ulogic;
    -- output
  );
end RSA_Core;
  
  
  
architecture behaviour of RSA_Core is
  -- internal signals
begin -- logic

end behaviour;
