

entity RSA is
  port(
    -- input
    -- output
  );
end RSA;
  
  
  
architecture behaviour of RSA is
  --internal signals
begin -- logic

end behaviour;
